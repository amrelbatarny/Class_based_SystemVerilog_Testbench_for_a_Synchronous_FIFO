package shared_pkg;
	int correct_count, error_count;
	bit test_finished;
endpackage : shared_pkg